module max2_test1(input ina, inb, output out);


assign out = ina & inb;

endmodule 