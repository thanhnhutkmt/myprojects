module myAnd(in1, in2, out);

input in1;
input in2;
wire in1;
wire in2;

output out;
reg out = in1 & in2;


endmodule 